(** Basically, this file just puts together all of the StackFrame stuff
  * in one place, so that I could refactor StackFrame into multiple files
  * but not have to rename the module everywhere *)

Require Export StackFrame1 StackFrameMinHelpers StackFrameMin.
